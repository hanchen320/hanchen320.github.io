-- amuntitled_GN.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity amuntitled_GN is
	port (
		SinDelay  : out std_logic_vector(15 downto 0);                    --  SinDelay.wire
		StreamMod : out std_logic_vector(18 downto 0);                    -- StreamMod.wire
		Noise     : in  std_logic                     := '0';             --     Noise.wire
		Sinln2    : out std_logic_vector(15 downto 0);                    --    Sinln2.wire
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		aclr      : in  std_logic                     := '0';             --          .reset
		Sinln     : in  std_logic_vector(15 downto 0) := (others => '0'); --     Sinln.wire
		StreamBit : out std_logic                                         -- StreamBit.wire
	);
end entity amuntitled_GN;

architecture rtl of amuntitled_GN is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_port_GN5RJOJIHL is
		port (
			input  : in  std_logic_vector(18 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(18 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GN5RJOJIHL;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_port_GNBO6OMO5Y is
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNBO6OMO5Y;

	component alt_dspbuilder_product_GNO6FDVQSR is
		generic (
			UseDedicatedMult : natural := 0;
			Signed           : natural := 0;
			lpm              : natural := 0;
			MaskValue        : string  := "1";
			pipeline         : natural := 0;
			width_b          : natural := 8;
			width_a          : natural := 8
		);
		port (
			aclr      : in  std_logic                                      := 'X';             -- clk
			clock     : in  std_logic                                      := 'X';             -- clk
			dataa     : in  std_logic_vector(width_a-1 downto 0)           := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width_b-1 downto 0)           := (others => 'X'); -- wire
			ena       : in  std_logic                                      := 'X';             -- wire
			result    : out std_logic_vector(width_a + width_b-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                      := 'X'              -- wire
		);
	end component alt_dspbuilder_product_GNO6FDVQSR;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_bus_build_GNGCK3JP43 is
		generic (
			width : natural := 8
		);
		port (
			output : out std_logic_vector(1 downto 0);        -- wire
			in0    : in  std_logic                    := 'X'; -- wire
			in1    : in  std_logic                    := 'X'  -- wire
		);
	end component alt_dspbuilder_bus_build_GNGCK3JP43;

	component alt_dspbuilder_delay_GNG36NZ2PG is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNG36NZ2PG;

	component alt_dspbuilder_cast_GN2TL7HGV4 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(1 downto 0) := (others => 'X'); -- wire
			output : out std_logic                                        -- wire
		);
	end component alt_dspbuilder_cast_GN2TL7HGV4;

	component alt_dspbuilder_cast_GNYH4N5SPJ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(18 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNYH4N5SPJ;

	signal productuser_aclrgnd_output_wire : std_logic;                     -- Productuser_aclrGND:output -> Product:user_aclr
	signal productenavcc_output_wire       : std_logic;                     -- ProductenaVCC:output -> Product:ena
	signal delaysclrgnd_output_wire        : std_logic;                     -- DelaysclrGND:output -> Delay:sclr
	signal delayenavcc_output_wire         : std_logic;                     -- DelayenaVCC:output -> Delay:ena
	signal gnd_output_wire                 : std_logic;                     -- GND:output -> Bus_Builder:in1
	signal noise_0_output_wire             : std_logic;                     -- Noise_0:output -> Bus_Builder:in0
	signal bus_builder_output_wire         : std_logic_vector(1 downto 0);  -- Bus_Builder:output -> [Product:datab, cast0:input]
	signal delay_output_wire               : std_logic_vector(15 downto 0); -- Delay:output -> SinDelay_0:input
	signal sinln_0_output_wire             : std_logic_vector(15 downto 0); -- Sinln_0:output -> [Delay:input, Product:dataa, Sinln2_0:input]
	signal cast0_output_wire               : std_logic;                     -- cast0:output -> StreamBit_0:input
	signal product_result_wire             : std_logic_vector(17 downto 0); -- Product:result -> cast1:input
	signal cast1_output_wire               : std_logic_vector(18 downto 0); -- cast1:output -> StreamMod_0:input
	signal clock_0_clock_output_clk        : std_logic;                     -- Clock_0:clock_out -> [Delay:clock, Product:clock]
	signal clock_0_clock_output_reset      : std_logic;                     -- Clock_0:aclr_out -> [Delay:aclr, Product:aclr]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	streammod_0 : component alt_dspbuilder_port_GN5RJOJIHL
		port map (
			input  => cast1_output_wire, --  input.wire
			output => StreamMod          -- output.wire
		);

	noise_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Noise,               --  input.wire
			output => noise_0_output_wire  -- output.wire
		);

	sinln2_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => sinln_0_output_wire, --  input.wire
			output => Sinln2               -- output.wire
		);

	product : component alt_dspbuilder_product_GNO6FDVQSR
		generic map (
			UseDedicatedMult => 1,
			Signed           => 1,
			lpm              => 0,
			MaskValue        => "1",
			pipeline         => 0,
			width_b          => 2,
			width_a          => 16
		)
		port map (
			clock     => clock_0_clock_output_clk,        -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,      --           .reset
			dataa     => sinln_0_output_wire,             --      dataa.wire
			datab     => bus_builder_output_wire,         --      datab.wire
			result    => product_result_wire,             --     result.wire
			user_aclr => productuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => productenavcc_output_wire        --        ena.wire
		);

	productuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => productuser_aclrgnd_output_wire  -- output.wire
		);

	productenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => productenavcc_output_wire  -- output.wire
		);

	bus_builder : component alt_dspbuilder_bus_build_GNGCK3JP43
		generic map (
			width => 2
		)
		port map (
			output => bus_builder_output_wire, -- output.wire
			in0    => noise_0_output_wire,     --    in0.wire
			in1    => gnd_output_wire          --    in1.wire
		);

	streambit_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => cast0_output_wire, --  input.wire
			output => StreamBit          -- output.wire
		);

	delay : component alt_dspbuilder_delay_GNG36NZ2PG
		generic map (
			ClockPhase => "1",
			BitPattern => "0000000000000001",
			width      => 16,
			use_init   => 0,
			delay      => 1
		)
		port map (
			input  => sinln_0_output_wire,        --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay_output_wire,          --     output.wire
			sclr   => delaysclrgnd_output_wire,   --       sclr.wire
			ena    => delayenavcc_output_wire     --        ena.wire
		);

	delaysclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delaysclrgnd_output_wire  -- output.wire
		);

	delayenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delayenavcc_output_wire  -- output.wire
		);

	sindelay_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => delay_output_wire, --  input.wire
			output => SinDelay           -- output.wire
		);

	sinln_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => Sinln,               --  input.wire
			output => sinln_0_output_wire  -- output.wire
		);

	gnd : component alt_dspbuilder_gnd_GN
		port map (
			output => gnd_output_wire  -- output.wire
		);

	cast0 : component alt_dspbuilder_cast_GN2TL7HGV4
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_builder_output_wire, --  input.wire
			output => cast0_output_wire        -- output.wire
		);

	cast1 : component alt_dspbuilder_cast_GNYH4N5SPJ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => product_result_wire, --  input.wire
			output => cast1_output_wire    -- output.wire
		);

end architecture rtl; -- of amuntitled_GN
