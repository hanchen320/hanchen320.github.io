-- tb_amuntitled.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb_amuntitled is
end entity tb_amuntitled;

architecture rtl of tb_amuntitled is
	component amuntitled_GN is
		port (
			Clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			StreamMod : out std_logic_vector(18 downto 0);                    -- wire
			Noise     : in  std_logic                     := 'X';             -- wire
			Sinln2    : out std_logic_vector(15 downto 0);                    -- wire
			StreamBit : out std_logic;                                        -- wire
			SinDelay  : out std_logic_vector(15 downto 0);                    -- wire
			Sinln     : in  std_logic_vector(15 downto 0) := (others => 'X')  -- wire
		);
	end component amuntitled_GN;

	component alt_dspbuilder_testbench_clock_GNCGUFKHRR is
		generic (
			SIMULATION_START_CYCLE       : natural := 4;
			RESET_REGISTER_CASCADE_DEPTH : natural := 0;
			RESET_LATENCY                : natural := 0
		);
		port (
			aclr_out     : out std_logic;  -- reset
			clock_out    : out std_logic;  -- clk
			reg_aclr_out : out std_logic;  -- reset
			tb_aclr      : out std_logic   -- reset
		);
	end component alt_dspbuilder_testbench_clock_GNCGUFKHRR;

	component alt_dspbuilder_testbench_salt_GNDBMPYDND is
		generic (
			XFILE : string := "default"
		);
		port (
			clock  : in  std_logic := 'X'; -- clk
			aclr   : in  std_logic := 'X'; -- reset
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_testbench_salt_GNDBMPYDND;

	component alt_dspbuilder_testbench_salt_GNQ2RNDGBK is
		generic (
			XFILE : string := "default"
		);
		port (
			clock  : in  std_logic                     := 'X'; -- clk
			aclr   : in  std_logic                     := 'X'; -- reset
			output : out std_logic_vector(15 downto 0)         -- wire
		);
	end component alt_dspbuilder_testbench_salt_GNQ2RNDGBK;

	component alt_dspbuilder_testbench_capture_GNUHQBGHYW is
		generic (
			DSPBTYPE : string := "";
			XFILE    : string := "default"
		);
		port (
			clock : in std_logic                     := 'X';             -- clk
			aclr  : in std_logic                     := 'X';             -- reset
			input : in std_logic_vector(18 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_testbench_capture_GNUHQBGHYW;

	component alt_dspbuilder_testbench_capture_GNAXODEVVW is
		generic (
			DSPBTYPE : string := "";
			XFILE    : string := "default"
		);
		port (
			clock : in std_logic                     := 'X';             -- clk
			aclr  : in std_logic                     := 'X';             -- reset
			input : in std_logic_vector(15 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_testbench_capture_GNAXODEVVW;

	component alt_dspbuilder_testbench_capture_GNQX2JTRTZ is
		generic (
			DSPBTYPE : string := "";
			XFILE    : string := "default"
		);
		port (
			clock : in std_logic := 'X'; -- clk
			aclr  : in std_logic := 'X'; -- reset
			input : in std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_testbench_capture_GNQX2JTRTZ;

	signal salt_noise_output_wire      : std_logic;                     -- salt_Noise:output -> dut:Noise
	signal clock_clock_tb_clk          : std_logic;                     -- Clock:clock_out -> [capture_SinDelay:clock, capture_Sinln2:clock, capture_StreamBit:clock, capture_StreamMod:clock, dut:Clock, salt_Noise:clock, salt_Sinln:clock]
	signal clock_clock_tb_reset        : std_logic;                     -- Clock:tb_aclr -> [salt_Noise:aclr, salt_Sinln:aclr]
	signal salt_sinln_output_wire      : std_logic_vector(15 downto 0); -- salt_Sinln:output -> dut:Sinln
	signal dut_streammod_wire          : std_logic_vector(18 downto 0); -- dut:StreamMod -> capture_StreamMod:input
	signal clock_clock_reg_reset_reset : std_logic;                     -- Clock:reg_aclr_out -> [capture_SinDelay:aclr, capture_Sinln2:aclr, capture_StreamBit:aclr, capture_StreamMod:aclr]
	signal dut_sinln2_wire             : std_logic_vector(15 downto 0); -- dut:Sinln2 -> capture_Sinln2:input
	signal dut_streambit_wire          : std_logic;                     -- dut:StreamBit -> capture_StreamBit:input
	signal dut_sindelay_wire           : std_logic_vector(15 downto 0); -- dut:SinDelay -> capture_SinDelay:input
	signal clock_clock_output_reset    : std_logic;                     -- Clock:aclr_out -> dut:aclr

begin

	dut : component amuntitled_GN
		port map (
			Clock     => clock_clock_tb_clk,       --     Clock.clk
			aclr      => clock_clock_output_reset, --          .reset
			StreamMod => dut_streammod_wire,       -- StreamMod.wire
			Noise     => salt_noise_output_wire,   --     Noise.wire
			Sinln2    => dut_sinln2_wire,          --    Sinln2.wire
			StreamBit => dut_streambit_wire,       -- StreamBit.wire
			SinDelay  => dut_sindelay_wire,        --  SinDelay.wire
			Sinln     => salt_sinln_output_wire    --     Sinln.wire
		);

	clock : component alt_dspbuilder_testbench_clock_GNCGUFKHRR
		generic map (
			SIMULATION_START_CYCLE       => 5,
			RESET_REGISTER_CASCADE_DEPTH => 0,
			RESET_LATENCY                => 0
		)
		port map (
			clock_out    => clock_clock_tb_clk,          --        clock_tb.clk
			tb_aclr      => clock_clock_tb_reset,        --                .reset
			aclr_out     => clock_clock_output_reset,    --    clock_output.reset
			reg_aclr_out => clock_clock_reg_reset_reset  -- clock_reg_reset.reset
		);

	salt_noise : component alt_dspbuilder_testbench_salt_GNDBMPYDND
		generic map (
			XFILE => "amuntitled_Noise.salt"
		)
		port map (
			clock  => clock_clock_tb_clk,     -- clock_aclr.clk
			aclr   => clock_clock_tb_reset,   --           .reset
			output => salt_noise_output_wire  --     output.wire
		);

	salt_sinln : component alt_dspbuilder_testbench_salt_GNQ2RNDGBK
		generic map (
			XFILE => "amuntitled_Sinln.salt"
		)
		port map (
			clock  => clock_clock_tb_clk,     -- clock_aclr.clk
			aclr   => clock_clock_tb_reset,   --           .reset
			output => salt_sinln_output_wire  --     output.wire
		);

	capture_streammod : component alt_dspbuilder_testbench_capture_GNUHQBGHYW
		generic map (
			DSPBTYPE => "INT [19, 0]",
			XFILE    => "amuntitled_StreamMod.capture.msim"
		)
		port map (
			clock => clock_clock_tb_clk,          -- clock_aclr.clk
			aclr  => clock_clock_reg_reset_reset, --           .reset
			input => dut_streammod_wire           --      input.wire
		);

	capture_sinln2 : component alt_dspbuilder_testbench_capture_GNAXODEVVW
		generic map (
			DSPBTYPE => "INT [16, 0]",
			XFILE    => "amuntitled_Sinln2.capture.msim"
		)
		port map (
			clock => clock_clock_tb_clk,          -- clock_aclr.clk
			aclr  => clock_clock_reg_reset_reset, --           .reset
			input => dut_sinln2_wire              --      input.wire
		);

	capture_streambit : component alt_dspbuilder_testbench_capture_GNQX2JTRTZ
		generic map (
			DSPBTYPE => "BIT [1, 0]",
			XFILE    => "amuntitled_StreamBit.capture.msim"
		)
		port map (
			clock => clock_clock_tb_clk,          -- clock_aclr.clk
			aclr  => clock_clock_reg_reset_reset, --           .reset
			input => dut_streambit_wire           --      input.wire
		);

	capture_sindelay : component alt_dspbuilder_testbench_capture_GNAXODEVVW
		generic map (
			DSPBTYPE => "INT [16, 0]",
			XFILE    => "amuntitled_SinDelay.capture.msim"
		)
		port map (
			clock => clock_clock_tb_clk,          -- clock_aclr.clk
			aclr  => clock_clock_reg_reset_reset, --           .reset
			input => dut_sindelay_wire            --      input.wire
		);

end architecture rtl; -- of tb_amuntitled
